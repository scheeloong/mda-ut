// RS232_0.v

// Generated using ACDS version 12.0 178 at 2012.09.26.10:29:14

`timescale 1 ps / 1 ps
module RS232_slave (
		input  wire        clk,        //            clock.clk
		input  wire        reset,      //            reset.reset
		input  wire        address,    //   avalon_slave_0.address
		input  wire        chipselect, //                 .chipselect
		input  wire [3:0]  byteenable, //                 .byteenable
		input  wire        read,       //                 .read
		input  wire        write,      //                 .write
		input  wire [31:0] writedata,  //                 .writedata
		output wire [31:0] readdata,   //                 .readdata
		input  wire        UART_RXD,   //      conduit_end.export
		output wire        UART_TXD,   //    conduit_end_1.export
		output wire        irq         // interrupt_sender.irq
	);

	Altera_UP_Avalon_RS232 rs232_0_inst (
		.clk        (clk),        //            clock.clk
		.reset      (reset),      //            reset.reset
		.address    (address),    //   avalon_slave_0.address
		.chipselect (chipselect), //                 .chipselect
		.byteenable (byteenable), //                 .byteenable
		.read       (read),       //                 .read
		.write      (write),      //                 .write
		.writedata  (writedata),  //                 .writedata
		.readdata   (readdata),   //                 .readdata
		.UART_RXD   (UART_RXD),   //      conduit_end.export
		.UART_TXD   (UART_TXD),   //    conduit_end_1.export
		.irq        (irq)         // interrupt_sender.irq
	);

endmodule
